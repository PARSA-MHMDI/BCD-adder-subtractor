library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity nines_compliment is
			port(
			
			);
end nines_compliment;

architecture Behavioral of nines_compliment is

begin


end Behavioral;

